
module soc_system (
	button_pio_external_connection_export,
	clk_clk,
	clk_freq_div_2_external_connection_export,
	dipsw_pio_external_connection_export,
	dispense_timer_external_connection_export,
	fisnar_inputs_external_connection_export,
	fisnar_outputs_external_connection_export,
	hps_0_f2h_cold_reset_req_reset_n,
	hps_0_f2h_debug_reset_req_reset_n,
	hps_0_f2h_stm_hw_events_stm_hwevents,
	hps_0_f2h_warm_reset_req_reset_n,
	hps_0_h2f_reset_reset_n,
	hps_0_hps_io_hps_io_emac1_inst_TX_CLK,
	hps_0_hps_io_hps_io_emac1_inst_TXD0,
	hps_0_hps_io_hps_io_emac1_inst_TXD1,
	hps_0_hps_io_hps_io_emac1_inst_TXD2,
	hps_0_hps_io_hps_io_emac1_inst_TXD3,
	hps_0_hps_io_hps_io_emac1_inst_RXD0,
	hps_0_hps_io_hps_io_emac1_inst_MDIO,
	hps_0_hps_io_hps_io_emac1_inst_MDC,
	hps_0_hps_io_hps_io_emac1_inst_RX_CTL,
	hps_0_hps_io_hps_io_emac1_inst_TX_CTL,
	hps_0_hps_io_hps_io_emac1_inst_RX_CLK,
	hps_0_hps_io_hps_io_emac1_inst_RXD1,
	hps_0_hps_io_hps_io_emac1_inst_RXD2,
	hps_0_hps_io_hps_io_emac1_inst_RXD3,
	hps_0_hps_io_hps_io_sdio_inst_CMD,
	hps_0_hps_io_hps_io_sdio_inst_D0,
	hps_0_hps_io_hps_io_sdio_inst_D1,
	hps_0_hps_io_hps_io_sdio_inst_CLK,
	hps_0_hps_io_hps_io_sdio_inst_D2,
	hps_0_hps_io_hps_io_sdio_inst_D3,
	hps_0_hps_io_hps_io_usb1_inst_D0,
	hps_0_hps_io_hps_io_usb1_inst_D1,
	hps_0_hps_io_hps_io_usb1_inst_D2,
	hps_0_hps_io_hps_io_usb1_inst_D3,
	hps_0_hps_io_hps_io_usb1_inst_D4,
	hps_0_hps_io_hps_io_usb1_inst_D5,
	hps_0_hps_io_hps_io_usb1_inst_D6,
	hps_0_hps_io_hps_io_usb1_inst_D7,
	hps_0_hps_io_hps_io_usb1_inst_CLK,
	hps_0_hps_io_hps_io_usb1_inst_STP,
	hps_0_hps_io_hps_io_usb1_inst_DIR,
	hps_0_hps_io_hps_io_usb1_inst_NXT,
	hps_0_hps_io_hps_io_spim1_inst_CLK,
	hps_0_hps_io_hps_io_spim1_inst_MOSI,
	hps_0_hps_io_hps_io_spim1_inst_MISO,
	hps_0_hps_io_hps_io_spim1_inst_SS0,
	hps_0_hps_io_hps_io_uart0_inst_RX,
	hps_0_hps_io_hps_io_uart0_inst_TX,
	hps_0_hps_io_hps_io_i2c0_inst_SDA,
	hps_0_hps_io_hps_io_i2c0_inst_SCL,
	hps_0_hps_io_hps_io_i2c1_inst_SDA,
	hps_0_hps_io_hps_io_i2c1_inst_SCL,
	hps_0_hps_io_hps_io_gpio_inst_GPIO09,
	hps_0_hps_io_hps_io_gpio_inst_GPIO35,
	hps_0_hps_io_hps_io_gpio_inst_GPIO40,
	hps_0_hps_io_hps_io_gpio_inst_GPIO53,
	hps_0_hps_io_hps_io_gpio_inst_GPIO54,
	hps_0_hps_io_hps_io_gpio_inst_GPIO61,
	joystick_external_connection_export,
	led_pio_external_connection_export,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	pololu_external_connection_export,
	reset_reset_n,
	teach_fpga2hps_external_connection_export,
	teach_hps2fpga_external_connection_export,
	x_motor_accelstep_pio_external_connection_export,
	x_motor_ctrl_pio_external_connection_export,
	x_motor_homeloc_pio_external_connection_export,
	x_motor_homespeed_pio_external_connection_export,
	x_motor_location_pio_external_connection_export,
	x_motor_lowerlimit_pio_external_connection_export,
	x_motor_max_speed_pio_external_connection_export,
	x_motor_min_speed_pio_external_connection_export,
	x_motor_status_pio_external_connection_export,
	x_motor_stepincrement_pio_external_connection_export,
	x_motor_target_pio_external_connection_export,
	x_motor_upperlimit_pio_external_connection_export,
	y_motor_accelstep_pio_external_connection_export,
	y_motor_ctrl_pio_external_connection_export,
	y_motor_homeloc_pio_external_connection_export,
	y_motor_homespeed_pio_external_connection_export,
	y_motor_location_pio_external_connection_export,
	y_motor_lowerlimit_pio_external_connection_export,
	y_motor_max_speed_pio_external_connection_export,
	y_motor_min_speed_pio_external_connection_export,
	y_motor_status_pio_external_connection_export,
	y_motor_stepincrement_pio_external_connection_export,
	y_motor_target_pio_external_connection_export,
	y_motor_upperlimit_pio_external_connection_export,
	z_motor_accelstep_pio_external_connection_export,
	z_motor_ctrl_pio_external_connection_export,
	z_motor_homeloc_pio_external_connection_export,
	z_motor_homespeed_pio_external_connection_export,
	z_motor_location_pio_external_connection_export,
	z_motor_lowerlimit_pio_external_connection_export,
	z_motor_max_speed_pio_external_connection_export,
	z_motor_min_speed_pio_external_connection_export,
	z_motor_status_pio_external_connection_export,
	z_motor_stepincrement_pio_external_connection_export,
	z_motor_target_pio_external_connection_export,
	z_motor_upperlimit_pio_external_connection_export);	

	input	[1:0]	button_pio_external_connection_export;
	input		clk_clk;
	output	[31:0]	clk_freq_div_2_external_connection_export;
	input	[3:0]	dipsw_pio_external_connection_export;
	output	[31:0]	dispense_timer_external_connection_export;
	input	[31:0]	fisnar_inputs_external_connection_export;
	output	[31:0]	fisnar_outputs_external_connection_export;
	input		hps_0_f2h_cold_reset_req_reset_n;
	input		hps_0_f2h_debug_reset_req_reset_n;
	input	[27:0]	hps_0_f2h_stm_hw_events_stm_hwevents;
	input		hps_0_f2h_warm_reset_req_reset_n;
	output		hps_0_h2f_reset_reset_n;
	output		hps_0_hps_io_hps_io_emac1_inst_TX_CLK;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD0;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD1;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD2;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD3;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD0;
	inout		hps_0_hps_io_hps_io_emac1_inst_MDIO;
	output		hps_0_hps_io_hps_io_emac1_inst_MDC;
	input		hps_0_hps_io_hps_io_emac1_inst_RX_CTL;
	output		hps_0_hps_io_hps_io_emac1_inst_TX_CTL;
	input		hps_0_hps_io_hps_io_emac1_inst_RX_CLK;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD1;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD2;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD3;
	inout		hps_0_hps_io_hps_io_sdio_inst_CMD;
	inout		hps_0_hps_io_hps_io_sdio_inst_D0;
	inout		hps_0_hps_io_hps_io_sdio_inst_D1;
	output		hps_0_hps_io_hps_io_sdio_inst_CLK;
	inout		hps_0_hps_io_hps_io_sdio_inst_D2;
	inout		hps_0_hps_io_hps_io_sdio_inst_D3;
	inout		hps_0_hps_io_hps_io_usb1_inst_D0;
	inout		hps_0_hps_io_hps_io_usb1_inst_D1;
	inout		hps_0_hps_io_hps_io_usb1_inst_D2;
	inout		hps_0_hps_io_hps_io_usb1_inst_D3;
	inout		hps_0_hps_io_hps_io_usb1_inst_D4;
	inout		hps_0_hps_io_hps_io_usb1_inst_D5;
	inout		hps_0_hps_io_hps_io_usb1_inst_D6;
	inout		hps_0_hps_io_hps_io_usb1_inst_D7;
	input		hps_0_hps_io_hps_io_usb1_inst_CLK;
	output		hps_0_hps_io_hps_io_usb1_inst_STP;
	input		hps_0_hps_io_hps_io_usb1_inst_DIR;
	input		hps_0_hps_io_hps_io_usb1_inst_NXT;
	output		hps_0_hps_io_hps_io_spim1_inst_CLK;
	output		hps_0_hps_io_hps_io_spim1_inst_MOSI;
	input		hps_0_hps_io_hps_io_spim1_inst_MISO;
	output		hps_0_hps_io_hps_io_spim1_inst_SS0;
	input		hps_0_hps_io_hps_io_uart0_inst_RX;
	output		hps_0_hps_io_hps_io_uart0_inst_TX;
	inout		hps_0_hps_io_hps_io_i2c0_inst_SDA;
	inout		hps_0_hps_io_hps_io_i2c0_inst_SCL;
	inout		hps_0_hps_io_hps_io_i2c1_inst_SDA;
	inout		hps_0_hps_io_hps_io_i2c1_inst_SCL;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO09;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO35;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO40;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO53;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO54;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO61;
	input	[31:0]	joystick_external_connection_export;
	output	[7:0]	led_pio_external_connection_export;
	output	[14:0]	memory_mem_a;
	output	[2:0]	memory_mem_ba;
	output		memory_mem_ck;
	output		memory_mem_ck_n;
	output		memory_mem_cke;
	output		memory_mem_cs_n;
	output		memory_mem_ras_n;
	output		memory_mem_cas_n;
	output		memory_mem_we_n;
	output		memory_mem_reset_n;
	inout	[31:0]	memory_mem_dq;
	inout	[3:0]	memory_mem_dqs;
	inout	[3:0]	memory_mem_dqs_n;
	output		memory_mem_odt;
	output	[3:0]	memory_mem_dm;
	input		memory_oct_rzqin;
	output	[31:0]	pololu_external_connection_export;
	input		reset_reset_n;
	input	[31:0]	teach_fpga2hps_external_connection_export;
	output	[31:0]	teach_hps2fpga_external_connection_export;
	output	[31:0]	x_motor_accelstep_pio_external_connection_export;
	output	[31:0]	x_motor_ctrl_pio_external_connection_export;
	output	[31:0]	x_motor_homeloc_pio_external_connection_export;
	output	[31:0]	x_motor_homespeed_pio_external_connection_export;
	input	[31:0]	x_motor_location_pio_external_connection_export;
	output	[31:0]	x_motor_lowerlimit_pio_external_connection_export;
	output	[31:0]	x_motor_max_speed_pio_external_connection_export;
	output	[31:0]	x_motor_min_speed_pio_external_connection_export;
	input	[31:0]	x_motor_status_pio_external_connection_export;
	output	[31:0]	x_motor_stepincrement_pio_external_connection_export;
	output	[31:0]	x_motor_target_pio_external_connection_export;
	output	[31:0]	x_motor_upperlimit_pio_external_connection_export;
	output	[31:0]	y_motor_accelstep_pio_external_connection_export;
	output	[31:0]	y_motor_ctrl_pio_external_connection_export;
	output	[31:0]	y_motor_homeloc_pio_external_connection_export;
	output	[31:0]	y_motor_homespeed_pio_external_connection_export;
	input	[31:0]	y_motor_location_pio_external_connection_export;
	output	[31:0]	y_motor_lowerlimit_pio_external_connection_export;
	output	[31:0]	y_motor_max_speed_pio_external_connection_export;
	output	[31:0]	y_motor_min_speed_pio_external_connection_export;
	input	[31:0]	y_motor_status_pio_external_connection_export;
	output	[31:0]	y_motor_stepincrement_pio_external_connection_export;
	output	[31:0]	y_motor_target_pio_external_connection_export;
	output	[31:0]	y_motor_upperlimit_pio_external_connection_export;
	output	[31:0]	z_motor_accelstep_pio_external_connection_export;
	output	[31:0]	z_motor_ctrl_pio_external_connection_export;
	output	[31:0]	z_motor_homeloc_pio_external_connection_export;
	output	[31:0]	z_motor_homespeed_pio_external_connection_export;
	input	[31:0]	z_motor_location_pio_external_connection_export;
	output	[31:0]	z_motor_lowerlimit_pio_external_connection_export;
	output	[31:0]	z_motor_max_speed_pio_external_connection_export;
	output	[31:0]	z_motor_min_speed_pio_external_connection_export;
	input	[31:0]	z_motor_status_pio_external_connection_export;
	output	[31:0]	z_motor_stepincrement_pio_external_connection_export;
	output	[31:0]	z_motor_target_pio_external_connection_export;
	output	[31:0]	z_motor_upperlimit_pio_external_connection_export;
endmodule
